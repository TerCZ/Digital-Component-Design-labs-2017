module pl_computer(resetn, clock, mem_clock, pc, inst, ealu, malu, walu, io_in, io_out);
// ?????? pipelined_computer??????????????? 1-1 ????????

    input  [12:0] io_in;
    output [44:0] io_out;
    // ??? IO

    input resetn, clock, mem_clock;
    // ??????? module ????????????????? resetn????? clock?
    // ????? clock ??????? mem_clock ???mem_clock ?????? ROM ?
    // ???? RAM ???????????????
    // ?????????????????????

    output [31:0] pc, inst, ealu, malu, walu;
    // ????????????????? wire ??

    wire [31:0] bpc, jpc, npc, pc4, ins, inst;
    // ??????????????????,?? 32 ?????IF ??????

    wire [31:0] dpc4, da, db, dimm;
    // ??????????????????,?? 32 ?????ID ???????

    wire [31:0] epc4, ea, eb, eimm;
    // ??????????????????,?? 32 ?????EXE ???????

    wire [31:0] mb, mmo;
    // ??????????????????,?? 32 ?????MEM ???????

    wire [31:0] wmo, wdi;
    // ??????????????????,?? 32 ?????WB ????????

    wire [4:0] drn, ern0, ern, mrn, wrn;
    // ????????????????????????????????32 ??? 5bit?

    wire [3:0] daluc, ealuc;
    // ID ??? EXE ????????????? aluc ?????4bit?

    wire [1:0] pcsource;
    // CU ??? IF ??????? PC ?????2bit?

    wire wpcir;
    // CU ??????????????????? PC ? IF/ID ???????????

    wire dwreg, dm2reg, dwmem, daluimm, dshift, djal;  // id stage
    // ID ??????????????????

    wire ewreg, em2reg, ewmem, ealuimm, eshift, ejal;  // exe stage
    // ??? ID/EXE ???????EXE ????????????????????

    wire mwreg, mm2reg, mwmem;  // mem stage
    // ??? EXE/MEM ???????MEM ????????????????????

    wire wwreg, wm2reg;  // wb stage
    // ??? MEM/WB ???????WB ????????

    pipepc prog_cnt(npc, wpcir, clock, resetn, pc);
    // ?????????????? IF ???????

    pipeif if_stage(pcsource, pc, bpc, da, jpc, npc, pc4, ins, mem_clock);  // IF stage
    // IF ????????????????? ROM ?????????
    // ???????? mem_clock ????????? rom_clk?
    // ???????? clock ??????? mem_clock??? rom_clock?,
    // ???????????????

    pipeir inst_reg(pc4, ins, wpcir, clock, resetn, dpc4, inst);  // IF/ID ??????
    // IF/ID ???????????? IF ??? ID ????????
    // ? clock ?????? IF ?????? ID ????????? IF/ID ??????
    // ?????? ID ???

    pipeid id_stage(mwreg, mrn, ern, ewreg, em2reg, mm2reg, dpc4, inst,
                    wrn, wdi, ealu, malu, mmo, wwreg, clock, resetn,
                    bpc, jpc, pcsource, wpcir, dwreg, dm2reg, dwmem, daluc,
                    daluimm, da, db, dimm, drn, dshift, djal);  // ID stage
    // ID ???????????????? CU??????????????
    // ???????????? clock ?????????????????? WB ??
    // ???????? clock ???????????????
    // ??? CU ???????????????????

    pipedereg de_reg(dwreg, dm2reg, dwmem, daluc, daluimm, da, db, dimm, drn, dshift,
                     djal, dpc4, clock, resetn, ewreg, em2reg, ewmem, ealuc, ealuimm,
                     ea, eb, eimm, ern0, eshift, ejal, epc4);  // ID/EXE ??????
    // ID/EXE ???????????? ID ??? EXE ????????
    // ? clock ?????? ID ?????? EXE ????????? ID/EXE ???
    // ????????? EXE ???

    pipeexe exe_stage(ealuc, ealuimm, ea, eb, eimm, eshift, ern0, epc4, ejal, ern, ealu);  // EXE stage
    // EXE ????????? ALU ????????

    pipeemreg em_reg(ewreg, em2reg, ewmem, ealu, eb, ern, clock, resetn,
                     mwreg, mm2reg, mwmem, malu, mb, mrn);  // EXE/MEM ??????
    // EXE/MEM ???????????? EXE ??? MEM ????????
    // ? clock ?????? EXE ?????? MEM ????????? EXE/MEM
    // ???????????? MEM ???

    pipemem mem_stage(mwmem, malu, mb, clock, mem_clock, mmo, io_in, io_out);  // MEM stage
    // MEM ???????????????? RAM ??????// ?? mem_clock?
    // ?????? RAM ? mem_clock ????????? ram_clk?
    // ???????? clock ??????? mem_clock ????? ram_clk?,
    // ?????????????????? mem_clock ?????????????

    pipemwreg mw_reg(mwreg, mm2reg, mmo, malu, mrn, clock, resetn,
                     wwreg, wm2reg, wmo, walu, wrn);  // MEM/WB ??????
    // MEM/WB ???????????? MEM ??? WB ????????
    // ? clock ?????? MEM ?????? WB ????????? MEM/WB
    // ???????????? WB ???

    mux2x32 wb_stage(walu, wmo, wm2reg, wdi);  // WB stage
    // WB ??????????????????????????????????
    // ??????????????????????????????
    // ?????????????????????
endmodule
